* SPICE3 file created from /home/raditya/Documents/Projects/Silicons/Projects/vco.ext - technology: sky130A

.option scale=10m

X0 a_1265_380# VCONT- a_985_380# VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X1 a_985_380# a_705_380# VGND VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X2 a_425_380# a_145_380# VGND VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X3 VGND a_705_380# sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X4 a_985_380# a_705_380# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X5 a_425_380# a_145_380# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X6 OUT a_1265_380# VGND VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X7 a_705_380# VCONT+ a_425_380# VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X8 a_145_380# VCONT+ OUT VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X9 VGND a_1265_380# sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X10 OUT a_1265_380# VPWR VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X11 a_705_380# VCONT- a_425_380# VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X12 VGND a_145_380# sky130_fd_pr__cap_mim_m3_1 l=1000 w=1000
X13 a_145_380# VCONT- OUT VPWR sky130_fd_pr__pfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
X14 a_1265_380# VCONT+ a_985_380# VGND sky130_fd_pr__nfet_01v8 ad=2.025n pd=0.18m as=2.025n ps=0.18m w=45 l=20
